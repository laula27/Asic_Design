// $Id: $
// File name:   tb_addernbit.sv
// Created:     2/3/2021
// Author:      Laula Student
// Lab Section: 337-015
// Version:     1.0  Initial Design Entry
// Description: postlab third
